/*
Cordic一次总旋转的前处理（预处理）：
将可能在4个象限任一象限中源向量[0°,360°) 映射到 第一象限的1/4象限中[0°, 45°)
*/
module cordic_pre(
	// 系统信号
	clk					,	// 时钟（clock）
	rst_n				,	// 复位（reset）
	
	// 一次Cordic总旋转前处理前的信号（源向量[0°,360°) ，故需要符号位）
	din_vsync			,	// 输入数据场有效信号
	din_hsync			,	// 输入数据行有效信号
	din_x				,	// 输入数据的x坐标（与 输入数据行有效信号 同步）
	din_y				,	// 输入数据的y坐标（与 输入数据行有效信号 同步）
	
	// 一次Cordic总旋转前处理后的信号（目的向量[0°, 45°)，故不需要符号位）
	dout_vsync			,	// 输出数据场有效信号
	dout_hsync			,	// 输出数据行有效信号
	dout_x				,	// 输出数据的x坐标（与 输出数据行有效信号 同步）
	dout_y				,	// 输出数据的y坐标（与 输出数据行有效信号 同步）
	// 输出源向量信息（与 输出数据行有效信号 同步）：
	// 第2位表示源向量x坐标符号（0表示正数，1表示负数），
	// 第1位表示源向量y坐标符号（0表示正数，1表示负数），
	// 第0位表示映射到第一象限后的x、y坐标是否需要经过互换才能继续映射到1/4象限（0表示不需要互换，1表示需要互换）。
	dout_info				// 输出源向量信息（与 输出数据行有效信号 同步）
	);
	
	
	// *******************************************参数声明***************************************
	// 视频数据流参数
	// 设x、y绝对值最大值为max_x_y，则最终迭代结果最大值不超过2*max_x_y，故需要保留一位用于迭代过程。
	// 即 输入数据x、y坐标的 最高位为符号位，次高位保留为0，
	// 即 输入数据x、y坐标的绝对值 保存在 低DW-2位
	parameter	DW			=	'd16		;	// 输入数据x、y坐标位宽
	// ******************************************************************************************
	
	
	// *******************************************端口声明***************************************
	// 系统信号
	input							clk					;	// 时钟（clock）
	input							rst_n				;	// 复位（reset）
	
	// 一次Cordic总旋转前处理前的信号（源向量[0°,360°) ，故需要符号位）
	input							din_vsync			;	// 输入数据场有效信号
	input							din_hsync			;	// 输入数据行有效信号
	input	signed	[DW-1:0]		din_x				;	// 输入数据的x坐标（与 输入数据行有效信号 同步）
	input	signed	[DW-1:0]		din_y				;	// 输入数据的y坐标（与 输入数据行有效信号 同步）
	
	// 一次Cordic总旋转前处理后的信号（目的向量[0°, 45°)，故不需要符号位）
	output							dout_vsync			;	// 输出数据场有效信号
	output							dout_hsync			;	// 输出数据行有效信号
	output	reg		[DW-1:0]		dout_x				;	// 输出数据的x坐标（与 输出数据行有效信号 同步）
	output	reg		[DW-1:0]		dout_y				;	// 输出数据的y坐标（与 输出数据行有效信号 同步）
	// 输出源向量信息（与 输出数据行有效信号 同步）：
	// 第2位表示源向量x坐标符号（0表示正数，1表示负数），
	// 第1位表示源向量y坐标符号（0表示正数，1表示负数），
	// 第0位表示映射到第一象限后的x、y坐标是否需要经过互换才能继续映射到1/4象限（0表示不需要互换，1表示需要互换）。
	output	reg		[ 2:0]			dout_info			;	// 输出源向量信息（与 输出数据行有效信号 同步）
	// *******************************************************************************************
	
	
	// *****************************************内部信号声明**************************************
	// 映射到第一象限中（即 x、y坐标都取绝对值）的信号
	reg			[DW-1:0]			x_abs				;	// 源x坐标的绝对值（源向量映射到第一象限后的x坐标）
	reg			[DW-1:0]			y_abs				;	// 源y坐标的绝对值（源向量映射到第一象限后的y坐标）
	reg								x_sign				;	// 源x坐标的符号（正数为0，负数为1）
	reg								y_sign				;	// 源y坐标的符号（正数为0，负数为1）
	
	// 映射到第一象限的1/4象限中（即 对于绝对值坐标：x<y时，x、y坐标互换；否则不变）的信号
	wire		[DW-1:0]			x_swap				;	// 绝对值x坐标的交换值（第一象限的向量映射到第一象限的1/4象限后的x坐标）
	wire		[DW-1:0]			y_swap				;	// 绝对值y坐标的交换值（第一象限的向量映射到第一象限的1/4象限后的y坐标）
	wire							is_swap				;	// 绝对值x坐标、绝对值y坐标 是否需要互换
	
	// 一次Cordic总旋转前处理前的 场、行同步信号 打拍
	reg								din_vsync_r0		;	// 输入数据场有效信号 打1拍
	reg								din_vsync_r1		;	// 输入数据场有效信号 打2拍
	reg								din_hsync_r0		;	// 输入数据行有效信号 打1拍
	reg								din_hsync_r1		;	// 输入数据行有效信号 打2拍
	// *******************************************************************************************
	
	
	// ---绝对值计算 函数---
	function [DW-1:0]abs;
		// 输入信号
		input	signed	[DW-1:0]	data_in	;	// 输入有符号数
		// 函数实现
		begin
			if(data_in[DW-1] == 1'b1) // 如果输入的有符号数最高位为1，则表明此输入为负数，故，要将负数的补码转化为正数的补码，则须将负数取反后+1
				abs = ~data_in + 1'b1;
			else // 如果输入的有符号数最高位为0，则表明此输入为正数，故，其绝对值为其本身
				abs = data_in;
		end
	endfunction
	// ------
	
	
	// ---将四个象限的源向量 映射到 第一象限中，并记录源向量的象限信息---
	// 即 求取源向量的x、y坐标的取绝对值，并记录源向量的x、y坐标的符号
	always @(posedge clk, negedge rst_n)
	begin
		if(!rst_n)
		begin
			x_abs <= 1'b0;
			y_abs <= 1'b0;
			x_sign <= 1'b0;
			y_sign <= 1'b0;
		end
		else if(din_hsync) // 输入有效时，开始转化、记录
		begin
			x_abs <= abs(din_x); // 调用绝对值函数 计算源x坐标的绝对值
			y_abs <= abs(din_y); // 调用绝对值函数 计算源y坐标的绝对值
			x_sign <= din_x[DW-1]; // 源有符号x坐标的最高位 记录了源x坐标的符号信息
			y_sign <= din_y[DW-1]; // 源有符号y坐标的最高位 记录了源y坐标的符号信息
		end
	end
	// ------
	
	
	// ---将第一象限的绝对值向量 映射到 第一象限的1/4象限中，并记录映射信息---
	// 即 对于绝对值坐标：当x<y时，x、y坐标互换；否则坐标不变。并记录是否互换了绝对值x、y坐标
	assign	is_swap	=	(x_abs<y_abs) ? 1'b1 : 1'b0	;
	assign	x_swap	=	is_swap ? y_abs : x_abs		;
	assign	y_swap	=	is_swap ? x_abs : y_abs		;
	// ------
	
	
	// ---最终映射到第一象限的1/4象限后的输出信号---
	// 最终映射到第一象限的1/4象限后的 x、y坐标，以及源向量信息
	always @(posedge clk, negedge rst_n)
	begin
		if(!rst_n)
		begin
			dout_x <= 1'b0;
			dout_y <= 1'b0;
			dout_info <= 1'b0;
		end
		else if(din_hsync_r0) // 有效期才输出
		begin
			dout_x <= x_swap;
			dout_y <= y_swap;
			dout_info <= {x_sign, y_sign, is_swap};
		end
		else
		begin
			dout_x <= 1'b0;
			dout_y <= 1'b0;
			dout_info <= 1'b0;
		end
	end
	
	// 一次Cordic总旋转前处理前的 场、行同步信号 打拍
	// 将四个象限的源向量 映射到 第一象限中，需要1个时钟；
	// 将第一象限的绝对值向量 映射到 第一象限的1/4象限中，需要1个时钟。
	// 即，从四个象限 映射到 第一象限的1/4象限，共需要2个时钟。
	// 故，场、行同步信号的输出也需要打2拍
	always @(posedge clk, negedge rst_n)
	begin
		if(!rst_n)
		begin
			din_vsync_r0 <= 1'b0;
			din_vsync_r1 <= 1'b0;
			din_hsync_r0 <= 1'b0;
			din_hsync_r1 <= 1'b0;
		end
		else
		begin
			din_vsync_r0 <= din_vsync;
			din_vsync_r1 <= din_vsync_r0;
			din_hsync_r0 <= din_hsync;
			din_hsync_r1 <= din_hsync_r0;
		end
	end
	
	// 最终映射到第一象限的1/4象限后的 场、行同步信号
	assign	dout_vsync	=	din_vsync_r1	;
	assign	dout_hsync	=	din_hsync_r1	;
	// ------
	
	
endmodule
