/*
Cordic一次总旋转（非伪旋转） 顶层模块：
将可能在4个象限任一象限中源向量[0°,360°) 经过一次Cordic总旋转，旋转到 0°轴上，
则旋转后的 x坐标即为 源向量的长度，y坐标即为 0，z坐标即为 源向量与0°轴的夹角的归一化值。
*/
module cordic_top(
	// 系统信号
	clk					,	// 时钟（clock）
	rst_n				,	// 复位（reset）
	
	// 一次Cordic总旋转前的信号（源向量[0°,360°) ，故需要符号位）
	din_vsync			,	// 输入数据场有效信号
	din_hsync			,	// 输入数据行有效信号
	din_x				,	// 输入数据的x坐标（与 输入数据行有效信号 同步）
	din_y				,	// 输入数据的y坐标（与 输入数据行有效信号 同步）
	
	// 一次Cordic总旋转后的信号（目的向量0°，故不需要符号位）
	dout_vsync			,	// 输出数据场有效信号
	dout_hsync			,	// 输出数据行有效信号
	dout_radians		,	// 输出源向量的模长（与 输出数据行有效信号 同步）
	dout_angle				// 输出源向量与0°轴的夹角α∈[0°, 360°)的归一化值：α/(2π)*(2^20)（与输出数据行有效信号同步）
	);
	
	
	// *******************************************参数声明***************************************
	// 视频数据流参数
	// 设x、y绝对值最大值为max_x_y，则最终迭代结果最大值不超过2*max_x_y，故需要保留一位用于迭代过程。
	// 即 输入数据x、y坐标的 最高位为符号位，次高位保留为0，
	// 即 输入数据x、y坐标的绝对值 保存在 低DW-2位
	parameter	DW			=	'd16		;	// 输入数据x、y坐标位宽
	
	// Cordic参数
	parameter	T_IR_NUM	=	'd15		;	// 总迭代次数（total iteration number）（可选 15~18）
	parameter	DW_DOT		=	'd4			;	// 输入数据x、y坐标的扩展小数位宽（用于提高精度）（输入数据x、y坐标位宽=DW+DW_DOT 须<=32）
	parameter	DW_NOR		=	'd20		;	// 输入数据z坐标归一化位宽（不要更改）
	// ******************************************************************************************
	
	
	// *******************************************端口声明***************************************
	// 系统信号
	input							clk					;	// 时钟（clock）
	input							rst_n				;	// 复位（reset）
	
	// 一次Cordic总旋转前的信号（源向量[0°,360°) ，故需要符号位）
	input							din_vsync			;	// 输入数据场有效信号
	input							din_hsync			;	// 输入数据行有效信号
	input	signed	[DW-1:0]		din_x				;	// 输入数据的x坐标（与 输入数据行有效信号 同步）
	input	signed	[DW-1:0]		din_y				;	// 输入数据的y坐标（与 输入数据行有效信号 同步）
	
	// 一次Cordic总旋转后的信号（目的向量0°，故不需要符号位）
	output							dout_vsync			;	// 输出数据场有效信号
	output							dout_hsync			;	// 输出数据行有效信号
	output			[DW-1:0]		dout_radians		;	// 输出源向量的模长（与 输出数据行有效信号 同步）
	output			[DW_NOR-1:0]	dout_angle			;	// 输出源向量与0°轴的夹角α∈[0°, 360°)的归一化值：α/(2π)*(2^20)（与输出数据行有效信号同步）
	// *******************************************************************************************
	
	
	// *****************************************内部信号声明**************************************
	// ---Cordic预处理模块信号---
	wire							pre_dout_vsync		;	// 预处理模块 输出数据场有效信号
	wire							pre_dout_hsync		;	// 预处理模块 输出数据行有效信号
	wire			[DW-1:0]		pre_dout_x			;	// 预处理模块 输出数据的x坐标（与 输出数据行有效信号 同步）
	wire			[DW-1:0]		pre_dout_y			;	// 预处理模块 输出数据的y坐标（与 输出数据行有效信号 同步）
	// 输出源向量信息（与 输出数据行有效信号 同步）：
	// 第2位表示源向量x坐标符号（0表示正数，1表示负数），
	// 第1位表示源向量y坐标符号（0表示正数，1表示负数），
	// 第0位表示映射到第一象限后的x、y坐标是否需要经过互换才能继续映射到1/4象限（0表示不需要互换，1表示需要互换）。
	wire			[ 2:0]			pre_dout_info		;	// 预处理模块 输出源向量信息（与 输出数据行有效信号 同步）
	
	// 预处理模块 输出源向量信息 打拍
	reg				[ 2:0]			pre_dout_info_r_arr[0:T_IR_NUM-1]	;	// 预处理模块输出源向量信息打T_IR_NUM拍
	// ------
	
	// ---Cordic总伪旋转模块信号---
	wire							core_dout_vsync		;	// 总伪旋转模块 输出数据场有效信号
	wire							core_dout_hsync		;	// 总伪旋转模块 输出数据行有效信号
	wire			[DW+DW_DOT-1:0]	core_dout_x			;	// 总伪旋转模块 输出数据的x坐标（与 输出数据行有效信号 同步）（扩展了小数位）
	wire			[DW_NOR-1:0]	core_dout_z			;	// 总伪旋转模块 输出数据的z坐标（与 输出数据行有效信号 同步）
	// ------
	
	// ---Cordic后处理模块信号---
	// 输入源向量信息（与 后处理输入数据行有效信号 同步）：
	// 第2位表示源向量x坐标符号（0表示正数，1表示负数），
	// 第1位表示源向量y坐标符号（0表示正数，1表示负数），
	// 第0位表示映射到第一象限后的x、y坐标是否需要经过互换才能继续映射到1/4象限（0表示不需要互换，1表示需要互换）。
	wire			[ 2:0]			post_din_info		;	// 后处理模块 输入源向量信息（与 后处理输入数据行有效信号 同步）
	// ------
	
	// for循环参数
	integer							i					;	// for循环计数值
	// *******************************************************************************************
	
	
	// ---实例化 Cordic一次总旋转的前处理（预处理） 模块---
	cordic_pre #(
		// 视频数据流参数
		// 设x、y绝对值最大值为max_x_y，则最终迭代结果最大值不超过2*max_x_y，故需要保留一位用于迭代过程。
		// 即 输入数据x、y坐标的 最高位为符号位，次高位保留为0，
		// 即 输入数据x、y坐标的绝对值 保存在 低DW-2位
		.DW					(DW				)	// 输入数据x、y坐标位宽
		)
	cordic_pre_u0(
		// 系统信号
		.clk				(clk			),	// 时钟（clock）
		.rst_n				(rst_n			),	// 复位（reset）
		
		// 一次Cordic总旋转前处理前的信号（源向量[0°,360°) ，故需要符号位）
		.din_vsync			(din_vsync		),	// 输入数据场有效信号
		.din_hsync			(din_hsync		),	// 输入数据行有效信号
		.din_x				(din_x			),	// 输入数据的x坐标（与 输入数据行有效信号 同步）
		.din_y				(din_y			),	// 输入数据的y坐标（与 输入数据行有效信号 同步）
		
		// 一次Cordic总旋转前处理后的信号（目的向量[0°, 45°)，故不需要符号位）
		.dout_vsync			(pre_dout_vsync	),	// 输出数据场有效信号
		.dout_hsync			(pre_dout_hsync	),	// 输出数据行有效信号
		.dout_x				(pre_dout_x		),	// 输出数据的x坐标（与 输出数据行有效信号 同步）
		.dout_y				(pre_dout_y		),	// 输出数据的y坐标（与 输出数据行有效信号 同步）
		// 输出源向量信息（与 输出数据行有效信号 同步）：
		// 第2位表示源向量x坐标符号（0表示正数，1表示负数），
		// 第1位表示源向量y坐标符号（0表示正数，1表示负数），
		// 第0位表示映射到第一象限后的x、y坐标是否需要经过互换才能继续映射到1/4象限（0表示不需要互换，1表示需要互换），
		.dout_info			(pre_dout_info	)	// 输出源向量信息（与 输出数据行有效信号 同步）
		);
	// ------
	
	
	// ---实例化 Cordic一次总旋转（伪旋转，未进行模长补偿） 模块---
	cordic_core #(
		// 视频数据流参数
		// 设x、y绝对值最大值为max_x_y，则最终迭代结果最大值不超过2*max_x_y，故需要保留一位用于迭代过程。
		// 即 输入数据x、y坐标的 最高位为符号位，次高位保留为0，
		// 即 输入数据x、y坐标的绝对值 保存在 低DW-2位
		.DW					(DW				),	// 输入数据x、y坐标位宽
		
		// Cordic参数
		.T_IR_NUM			(T_IR_NUM		),	// 总迭代次数（total iteration number）（可选 15~18）
		.DW_DOT				(DW_DOT			)	// 输入数据x、y坐标的扩展小数位宽（用于提高精度）（输出数据x、y坐标位宽=DW+DW_DOT 须<=32）
		)
	cordic_core_u0(
		// 系统信号
		.clk				(clk			),	// 时钟（clock）
		.rst_n				(rst_n			),	// 复位（reset）
		
		// 一次Cordic总旋转前的信号
		// （因为是从0°~45°位置开始旋转的，也就是第一象限的1/4象限，故开始旋转前，x、y均>=0，而z取方向为从0到目标角 即 z=0，故x、y、z均不需要有符号位）
		.din_vsync			(pre_dout_vsync	),	// 输入数据场有效信号
		.din_hsync			(pre_dout_hsync	),	// 输入数据行有效信号
		.din_x				(pre_dout_x		),	// 输入数据的x坐标（与 输入数据行有效信号 同步）
		.din_y				(pre_dout_y		),	// 输入数据的y坐标（与 输入数据行有效信号 同步）
		.din_z				({DW_NOR{1'b0}}	),	// 输入数据的z坐标（与 输入数据行有效信号 同步）
		
		// 一次Cordic总旋转后的信号
		// （因为最终旋转到0°，故总旋转后，x>0，y坐标一定趋近于0 即 不需要输出y坐标，
		// 而起始总旋转位置为第一象限的1/4象限，故总旋转后，z趋近于起始旋转角度 即 z>=0，故x、z均不需要符号位）
		.dout_vsync			(core_dout_vsync),	// 输出数据场有效信号
		.dout_hsync			(core_dout_hsync),	// 输出数据行有效信号
		.dout_x				(core_dout_x	),	// 输出数据的x坐标（与 输出数据行有效信号 同步）
		.dout_z				(core_dout_z	)	// 输出数据的z坐标（与 输出数据行有效信号 同步）
		);
	// ------
	
	
	// ---实例化 Cordic一次总旋转（伪旋转）的后处理 模块---
	cordic_post #(
		// 视频数据流参数
		.DW					(DW				),	// 输出数据x、y坐标位宽
		
		// Cordic参数
		.T_IR_NUM			(T_IR_NUM		),	// 总迭代次数（total iteration number）（可选 15~18）
		.DW_DOT				(DW_DOT			)	// 输入数据x、y坐标的扩展小数位宽（用于提高精度）（输入数据x、y坐标位宽=DW+DW_DOT 须<=32）
		)
	cordic_post_u0(
		// 系统信号
		.clk				(clk			),	// 时钟（clock）
		.rst_n				(rst_n			),	// 复位（reset）
		
		// 一次Cordic总旋转（伪旋转）后处理前的信号
		.din_vsync			(core_dout_vsync),	// 输入数据场有效信号
		.din_hsync			(core_dout_hsync),	// 输入数据行有效信号
		.din_x				(core_dout_x	),	// 输入数据的x坐标（与 输入数据行有效信号 同步）
		.din_z				(core_dout_z	),	// 输入数据的z坐标（与 输入数据行有效信号 同步）
		// 输入总旋转前的源向量信息（与 输出数据行有效信号 同步）：
		// 第2位表示源向量x坐标符号（0表示正数，1表示负数），
		// 第1位表示源向量y坐标符号（0表示正数，1表示负数），
		// 第0位表示映射到第一象限后的x、y坐标是否需要经过互换才能继续映射到1/4象限（0表示不需要互换，1表示需要互换）。
		.din_info			(post_din_info	),	// 输入总旋转前的源向量信息（与 输出数据行有效信号 同步）
		
		// 一次Cordic总旋转（伪旋转）后处理后的信号
		.dout_vsync			(dout_vsync		),	// 输出数据场有效信号
		.dout_hsync			(dout_hsync		),	// 输出数据行有效信号
		.dout_x				(dout_radians	),	// 输出数据的x坐标（与 输出数据行有效信号 同步）（源向量的模长）
		.dout_z				(dout_angle		)	// 输出数据的z坐标（源向量与0°轴的夹角α∈[0°, 360°)的归一化值：α/(2π)*(2^20)）
		);
	// 预处理模块 输出源向量信息 打T_IR_NUM拍
	// 因为预处理模块输出后，又经过了总伪旋转模块，才来到后处理模块，
	// 而总伪旋转模块的输出比其输入滞后了T_IR_NUM拍，
	// 所以 对于从预处理模块输出的源向量象限信号，若要作为后处理模块输入，则需要打T_IR_NUM拍
	always @(posedge clk, negedge rst_n)
	begin
		if(!rst_n)
		begin
			for(i=0; i<T_IR_NUM; i=i+1)
				pre_dout_info_r_arr[i] <= 1'b0;
		end
		else
		begin
			pre_dout_info_r_arr[0] <= pre_dout_info;
			for(i=1; i<T_IR_NUM; i=i+1)
				pre_dout_info_r_arr[i] <= pre_dout_info_r_arr[i-1];
		end
	end
	assign	post_din_info	=	pre_dout_info_r_arr[T_IR_NUM-1];
	// ------
	
	
endmodule
